library verilog;
use verilog.vl_types.all;
entity controller is
    generic(
        ir_fetch        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        decode          : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        ALU             : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        Reg_write       : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        ADI             : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        ADI_w           : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        LW1             : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        LW2             : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        SW2             : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        BEQ1            : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        BEQ2            : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        JLR1            : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        JLR2            : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi0);
        LHI             : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi1);
        JAL2            : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi0);
        Counter         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        LM1             : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        LM2             : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi1);
        SM1             : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi0);
        SM2             : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi1);
        SM3             : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi0);
        \Reset\         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi1)
    );
    port(
        clk             : in     vl_logic;
        count           : in     vl_logic_vector(3 downto 0);
        enable          : out    vl_logic;
        reset           : out    vl_logic;
        reset_pin       : in     vl_logic;
        load            : out    vl_logic;
        op_sel          : out    vl_logic_vector(1 downto 0);
        regw            : out    vl_logic;
        rw              : out    vl_logic_vector(1 downto 0);
        mux_ccr_sel     : out    vl_logic;
        mux_memw_sel    : out    vl_logic;
        mux_a_sel       : out    vl_logic_vector(1 downto 0);
        mux_B_sel       : out    vl_logic;
        mux_adi_sel     : out    vl_logic;
        mux_alu_sel     : out    vl_logic_vector(1 downto 0);
        mux_mem_sel     : out    vl_logic;
        mux_reg_sel     : out    vl_logic_vector(1 downto 0);
        mux_pc_sel      : out    vl_logic_vector(1 downto 0);
        mux_pcw_sel     : out    vl_logic_vector(1 downto 0);
        opcode          : in     vl_logic_vector(15 downto 0);
        cz              : in     vl_logic_vector(1 downto 0);
        wa              : out    vl_logic;
        wb              : out    vl_logic;
        wmdr            : out    vl_logic;
        wccr            : out    vl_logic;
        walu            : out    vl_logic;
        wir             : out    vl_logic;
        equal           : in     vl_logic;
        aorb            : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ir_fetch : constant is 1;
    attribute mti_svvh_generic_type of decode : constant is 1;
    attribute mti_svvh_generic_type of ALU : constant is 1;
    attribute mti_svvh_generic_type of Reg_write : constant is 1;
    attribute mti_svvh_generic_type of ADI : constant is 1;
    attribute mti_svvh_generic_type of ADI_w : constant is 1;
    attribute mti_svvh_generic_type of LW1 : constant is 1;
    attribute mti_svvh_generic_type of LW2 : constant is 1;
    attribute mti_svvh_generic_type of SW2 : constant is 1;
    attribute mti_svvh_generic_type of BEQ1 : constant is 1;
    attribute mti_svvh_generic_type of BEQ2 : constant is 1;
    attribute mti_svvh_generic_type of JLR1 : constant is 1;
    attribute mti_svvh_generic_type of JLR2 : constant is 1;
    attribute mti_svvh_generic_type of LHI : constant is 1;
    attribute mti_svvh_generic_type of JAL2 : constant is 1;
    attribute mti_svvh_generic_type of Counter : constant is 1;
    attribute mti_svvh_generic_type of LM1 : constant is 1;
    attribute mti_svvh_generic_type of LM2 : constant is 1;
    attribute mti_svvh_generic_type of SM1 : constant is 1;
    attribute mti_svvh_generic_type of SM2 : constant is 1;
    attribute mti_svvh_generic_type of SM3 : constant is 1;
    attribute mti_svvh_generic_type of \Reset\ : constant is 1;
end controller;
