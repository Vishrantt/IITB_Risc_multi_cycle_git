module memory(data_in,data_outs,addr,clk,rw);

input [15:0] data_in;
input clk;
input [1:0] rw;
input [5:0] addr;

reg [15:0] Memory [64:0];

output [15:0] data_outs;
reg [15:0] data_outs;


initial 
begin										
//Memory[0] <= 16'b0000_000_111_010_0_00;//  ADD									
//Memory[0] <= 16'b0000_000_010_000_0_10;//  ADC									
//Memory[0] <= 16'b0000_000_010_000_0_01;//  ADZ									
//Memory[0] <= 16'b0010_000_010_000_0_00;//  NDU									
//Memory[0] <= 16'b0010_000_010_000_0_10;//  NDC									
//Memory[0] <= 16'b0010_000_010_000_0_01;//  NDZ				
//Memory[0] <= 16'b0001_000_010_000001;  //  ADI					
//Memory[0] <= 16'b0011_000_111000001;   //  LHI								
//Memory[0] <= 16'b0100_000_010_000010;  //  LW					
//Memory[0] <= 16'b0101_000_010_000010;  //  SW
//Memory[0] <= 16'b0110_000_0_01011011;  //	LM	
//Memory[0] <= 16'b0111_000_0_00110101;  //  SM				
//Memory[0] <= 16'b1100_000_010_000001;  //  BEQ	
//Memory[0] <= 16'b1000_000_010000001;   //  JAL	
//Memory[0] <= 16'b1001_000_010_000011;  //  JLR
				

//Memory[0] <= 16'b1000_000_00001_1100;  	
//Memory[1] <= 16'b0100100110000101;
//Memory[2] <= 16'b0100110110000101;	
//Memory[3] <= 16'b0100000101010100;
//Memory[4] <= 16'b0100001101010101;
//Memory[5] <= 16'b0001000010000000;
//Memory[6] <= 16'b0010000001011000;
//Memory[7] <= 16'b0010011011011000;
//Memory[8] <= 16'b0001011011000000;
//Memory[9] <= 16'b0000100010100001;
//Memory[10] <= 16'b0000000000000000;
//Memory[11] <= 16'b0010110110110010;
//Memory[12] <= 16'b1100110101111010;
//Memory[13] <= 16'b0101100101010110;
//Memory[20] <= 16'h0001;
//Memory[21] <= 16'h000F;
//Memory[22] <= 16'h000C;
//Memory[23] <= 16'h0015;
//Memory[24] <= 16'h0003;
//Memory[25] <= 16'h0000;
//Memory[26] <= 16'h0045;
//Memory[29] <= 16'b0001011011000001;
//Memory[30] <= 16'b0001110110010111;
//Memory[31] <= 16'b0101000110000100;
//Memory[32] <= 16'b0100000110000000;
//Memory[33] <= 16'b0100001110000001;
//Memory[34] <= 16'b1100101001001011;
//Memory[35] <= 16'b0000000010010000;
//Memory[36] <= 16'b0000011100100010;
//Memory[37] <= 16'b0001001001111111;
//Memory[38] <= 16'b0001111111111011;
//
//Memory[46] <= 16'b0101010110000010;
//Memory[47] <= 16'b0101100110000011;
//Memory[48] <= 16'b0001011011111111;
//Memory[49] <= 16'b0101011110000101;
//Memory[50] <= 16'b0100111110000100;   Without LMSM

//with LM and SM				
//From 0 to 13

Memory[0] <= 16'b1000000000011100;
Memory[1] <= 16'b0100100110000101;
Memory[2] <= 16'b0001110000111101;
Memory[3] <= 16'b0100110110000101;
Memory[4] <= 16'b0110_000_000000011;

Memory[5] <= 16'b0001000010000000;
Memory[6] <= 16'b0010000001011000;
Memory[7] <= 16'b0010011011011000;
Memory[8] <= 16'b0001011011000000;
Memory[9] <= 16'b0000100010100001;
Memory[10] <= 16'b0000000000000000;
Memory[11] <= 16'b0010110110110010;
Memory[12] <= 16'b110011010111_1001;
Memory[13] <= 16'b0101100101010110;

//From 20 to 27
//Memory[20] <= 16'h0001;
//Memory[21] <= 16'h000F;
//Memory[22] <= 16'h000C;
//Memory[23] <= 16'hFFFF;
//Memory[24] <= 16'h0045;
//Memory[25] <= 16'hFFBB;
//Memory[26] <= 16'h0000;
//Memory[27] <= 16'h0000;
Memory[20] <= 16'h0001;
Memory[21] <= 16'h000F;
Memory[22] <= 16'h0000;
Memory[23] <= 16'h0015;
Memory[24] <= 16'h0003;
Memory[25] <= 16'h0000;
Memory[26] <= 16'h0045;

//From 29 to 38;
Memory[29] <= 16'b0001011011000001;
Memory[30] <= 16'b0001110110010111;
Memory[31] <= 16'b0101000110000100;
Memory[32] <= 16'b0100000110000000;
Memory[33] <= 16'b0100001110000001;
Memory[34] <= 16'b1100101001001011;
Memory[35] <= 16'b0000000010010000;
Memory[36] <= 16'b0000011100100010;
Memory[37] <= 16'b0001001001111111;
Memory[38] <= 16'b0001111111111011;

//From 46 to 50
Memory[46] <= 16'b0001110000000010;
Memory[47] <= 16'b0111_000_0_00010100;
Memory[48] <= 16'b0001011011111111;
Memory[49] <= 16'b0101011110000101;
Memory[50] <= 16'b0100111110000100;

end


always @ (posedge clk)
begin
	if (rw == 2'b01)
	Memory[addr] <= data_in;	
end

always @ (*)
begin 
	if (rw == 2'b10)
	data_outs <= Memory[addr];
	else
	data_outs <= 16'b0;
end

endmodule
